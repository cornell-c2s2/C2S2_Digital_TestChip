magic
tech sky130A
magscale 1 2
timestamp 1685998435
<< obsli1 >>
rect 1104 2159 462852 581553
<< obsm1 >>
rect 934 2128 463114 583160
<< metal2 >>
rect 12990 583200 13046 584000
rect 38750 583200 38806 584000
rect 64510 583200 64566 584000
rect 90270 583200 90326 584000
rect 116030 583200 116086 584000
rect 141790 583200 141846 584000
rect 167550 583200 167606 584000
rect 193310 583200 193366 584000
rect 219070 583200 219126 584000
rect 244830 583200 244886 584000
rect 270590 583200 270646 584000
rect 296350 583200 296406 584000
rect 322110 583200 322166 584000
rect 347870 583200 347926 584000
rect 373630 583200 373686 584000
rect 399390 583200 399446 584000
rect 425150 583200 425206 584000
rect 450910 583200 450966 584000
rect 115938 0 115994 800
rect 347870 0 347926 800
<< obsm2 >>
rect 938 583144 12934 583200
rect 13102 583144 38694 583200
rect 38862 583144 64454 583200
rect 64622 583144 90214 583200
rect 90382 583144 115974 583200
rect 116142 583144 141734 583200
rect 141902 583144 167494 583200
rect 167662 583144 193254 583200
rect 193422 583144 219014 583200
rect 219182 583144 244774 583200
rect 244942 583144 270534 583200
rect 270702 583144 296294 583200
rect 296462 583144 322054 583200
rect 322222 583144 347814 583200
rect 347982 583144 373574 583200
rect 373742 583144 399334 583200
rect 399502 583144 425094 583200
rect 425262 583144 450854 583200
rect 451022 583144 463110 583200
rect 938 856 463110 583144
rect 938 800 115882 856
rect 116050 800 347814 856
rect 347982 800 463110 856
<< metal3 >>
rect 463200 565224 464000 565344
rect 463200 528776 464000 528896
rect 463200 492328 464000 492448
rect 463200 455880 464000 456000
rect 0 437928 800 438048
rect 463200 419432 464000 419552
rect 463200 382984 464000 383104
rect 463200 346536 464000 346656
rect 463200 310088 464000 310208
rect 463200 273640 464000 273760
rect 463200 237192 464000 237312
rect 463200 200744 464000 200864
rect 463200 164296 464000 164416
rect 0 145936 800 146056
rect 463200 127848 464000 127968
rect 463200 91400 464000 91520
rect 463200 54952 464000 55072
rect 463200 18504 464000 18624
<< obsm3 >>
rect 800 565424 463200 581569
rect 800 565144 463120 565424
rect 800 528976 463200 565144
rect 800 528696 463120 528976
rect 800 492528 463200 528696
rect 800 492248 463120 492528
rect 800 456080 463200 492248
rect 800 455800 463120 456080
rect 800 438128 463200 455800
rect 880 437848 463200 438128
rect 800 419632 463200 437848
rect 800 419352 463120 419632
rect 800 383184 463200 419352
rect 800 382904 463120 383184
rect 800 346736 463200 382904
rect 800 346456 463120 346736
rect 800 310288 463200 346456
rect 800 310008 463120 310288
rect 800 273840 463200 310008
rect 800 273560 463120 273840
rect 800 237392 463200 273560
rect 800 237112 463120 237392
rect 800 200944 463200 237112
rect 800 200664 463120 200944
rect 800 164496 463200 200664
rect 800 164216 463120 164496
rect 800 146136 463200 164216
rect 880 145856 463200 146136
rect 800 128048 463200 145856
rect 800 127768 463120 128048
rect 800 91600 463200 127768
rect 800 91320 463120 91600
rect 800 55152 463200 91320
rect 800 54872 463120 55152
rect 800 18704 463200 54872
rect 800 18424 463120 18704
rect 800 2143 463200 18424
<< metal4 >>
rect 4208 2128 4528 581584
rect 19568 2128 19888 581584
rect 34928 2128 35248 581584
rect 50288 2128 50608 581584
rect 65648 2128 65968 581584
rect 81008 2128 81328 581584
rect 96368 2128 96688 581584
rect 111728 2128 112048 581584
rect 127088 2128 127408 581584
rect 142448 2128 142768 581584
rect 157808 2128 158128 581584
rect 173168 2128 173488 581584
rect 188528 2128 188848 581584
rect 203888 2128 204208 581584
rect 219248 2128 219568 581584
rect 234608 2128 234928 581584
rect 249968 2128 250288 581584
rect 265328 2128 265648 581584
rect 280688 2128 281008 581584
rect 296048 2128 296368 581584
rect 311408 2128 311728 581584
rect 326768 2128 327088 581584
rect 342128 2128 342448 581584
rect 357488 2128 357808 581584
rect 372848 2128 373168 581584
rect 388208 2128 388528 581584
rect 403568 2128 403888 581584
rect 418928 2128 419248 581584
rect 434288 2128 434608 581584
rect 449648 2128 449968 581584
<< obsm4 >>
rect 70163 4931 80928 581229
rect 81408 4931 96288 581229
rect 96768 4931 111648 581229
rect 112128 4931 127008 581229
rect 127488 4931 142368 581229
rect 142848 4931 157728 581229
rect 158208 4931 173088 581229
rect 173568 4931 188448 581229
rect 188928 4931 203808 581229
rect 204288 4931 219168 581229
rect 219648 4931 234528 581229
rect 235008 4931 249888 581229
rect 250368 4931 265248 581229
rect 265728 4931 280608 581229
rect 281088 4931 295968 581229
rect 296448 4931 311328 581229
rect 311808 4931 326688 581229
rect 327168 4931 342048 581229
rect 342528 4931 357408 581229
rect 357888 4931 372768 581229
rect 373248 4931 388128 581229
rect 388608 4931 403488 581229
rect 403968 4931 406029 581229
<< labels >>
rlabel metal3 s 463200 18504 464000 18624 6 adapter_parity
port 1 nsew signal output
rlabel metal2 s 115938 0 115994 800 6 clk
port 2 nsew signal input
rlabel metal3 s 463200 54952 464000 55072 6 io_oeb[0]
port 3 nsew signal output
rlabel metal2 s 322110 583200 322166 584000 6 io_oeb[10]
port 4 nsew signal output
rlabel metal2 s 270590 583200 270646 584000 6 io_oeb[11]
port 5 nsew signal output
rlabel metal2 s 219070 583200 219126 584000 6 io_oeb[12]
port 6 nsew signal output
rlabel metal2 s 167550 583200 167606 584000 6 io_oeb[13]
port 7 nsew signal output
rlabel metal2 s 116030 583200 116086 584000 6 io_oeb[14]
port 8 nsew signal output
rlabel metal2 s 64510 583200 64566 584000 6 io_oeb[15]
port 9 nsew signal output
rlabel metal2 s 12990 583200 13046 584000 6 io_oeb[16]
port 10 nsew signal output
rlabel metal3 s 0 145936 800 146056 6 io_oeb[17]
port 11 nsew signal output
rlabel metal3 s 463200 127848 464000 127968 6 io_oeb[1]
port 12 nsew signal output
rlabel metal3 s 463200 200744 464000 200864 6 io_oeb[2]
port 13 nsew signal output
rlabel metal3 s 463200 273640 464000 273760 6 io_oeb[3]
port 14 nsew signal output
rlabel metal3 s 463200 346536 464000 346656 6 io_oeb[4]
port 15 nsew signal output
rlabel metal3 s 463200 419432 464000 419552 6 io_oeb[5]
port 16 nsew signal output
rlabel metal3 s 463200 492328 464000 492448 6 io_oeb[6]
port 17 nsew signal output
rlabel metal3 s 463200 565224 464000 565344 6 io_oeb[7]
port 18 nsew signal output
rlabel metal2 s 425150 583200 425206 584000 6 io_oeb[8]
port 19 nsew signal output
rlabel metal2 s 373630 583200 373686 584000 6 io_oeb[9]
port 20 nsew signal output
rlabel metal2 s 141790 583200 141846 584000 6 master_cs
port 21 nsew signal output
rlabel metal2 s 90270 583200 90326 584000 6 master_miso
port 22 nsew signal input
rlabel metal2 s 38750 583200 38806 584000 6 master_mosi
port 23 nsew signal output
rlabel metal3 s 0 437928 800 438048 6 master_sclk
port 24 nsew signal output
rlabel metal3 s 463200 164296 464000 164416 6 minion_cs
port 25 nsew signal input
rlabel metal3 s 463200 455880 464000 456000 6 minion_cs_2
port 26 nsew signal input
rlabel metal2 s 347870 583200 347926 584000 6 minion_cs_3
port 27 nsew signal input
rlabel metal3 s 463200 382984 464000 383104 6 minion_miso
port 28 nsew signal output
rlabel metal2 s 399390 583200 399446 584000 6 minion_miso_2
port 29 nsew signal output
rlabel metal2 s 193310 583200 193366 584000 6 minion_miso_3
port 30 nsew signal output
rlabel metal3 s 463200 237192 464000 237312 6 minion_mosi
port 31 nsew signal input
rlabel metal3 s 463200 528776 464000 528896 6 minion_mosi_2
port 32 nsew signal input
rlabel metal2 s 296350 583200 296406 584000 6 minion_mosi_3
port 33 nsew signal input
rlabel metal3 s 463200 91400 464000 91520 6 minion_parity
port 34 nsew signal output
rlabel metal3 s 463200 310088 464000 310208 6 minion_sclk
port 35 nsew signal input
rlabel metal2 s 450910 583200 450966 584000 6 minion_sclk_2
port 36 nsew signal input
rlabel metal2 s 244830 583200 244886 584000 6 minion_sclk_3
port 37 nsew signal input
rlabel metal2 s 347870 0 347926 800 6 reset
port 38 nsew signal input
rlabel metal4 s 4208 2128 4528 581584 6 vccd1
port 39 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 581584 6 vccd1
port 39 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 581584 6 vccd1
port 39 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 581584 6 vccd1
port 39 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 581584 6 vccd1
port 39 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 581584 6 vccd1
port 39 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 581584 6 vccd1
port 39 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 581584 6 vccd1
port 39 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 581584 6 vccd1
port 39 nsew power bidirectional
rlabel metal4 s 280688 2128 281008 581584 6 vccd1
port 39 nsew power bidirectional
rlabel metal4 s 311408 2128 311728 581584 6 vccd1
port 39 nsew power bidirectional
rlabel metal4 s 342128 2128 342448 581584 6 vccd1
port 39 nsew power bidirectional
rlabel metal4 s 372848 2128 373168 581584 6 vccd1
port 39 nsew power bidirectional
rlabel metal4 s 403568 2128 403888 581584 6 vccd1
port 39 nsew power bidirectional
rlabel metal4 s 434288 2128 434608 581584 6 vccd1
port 39 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 581584 6 vssd1
port 40 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 581584 6 vssd1
port 40 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 581584 6 vssd1
port 40 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 581584 6 vssd1
port 40 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 581584 6 vssd1
port 40 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 581584 6 vssd1
port 40 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 581584 6 vssd1
port 40 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 581584 6 vssd1
port 40 nsew ground bidirectional
rlabel metal4 s 265328 2128 265648 581584 6 vssd1
port 40 nsew ground bidirectional
rlabel metal4 s 296048 2128 296368 581584 6 vssd1
port 40 nsew ground bidirectional
rlabel metal4 s 326768 2128 327088 581584 6 vssd1
port 40 nsew ground bidirectional
rlabel metal4 s 357488 2128 357808 581584 6 vssd1
port 40 nsew ground bidirectional
rlabel metal4 s 388208 2128 388528 581584 6 vssd1
port 40 nsew ground bidirectional
rlabel metal4 s 418928 2128 419248 581584 6 vssd1
port 40 nsew ground bidirectional
rlabel metal4 s 449648 2128 449968 581584 6 vssd1
port 40 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 464000 584000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 387920002
string GDS_FILE /home/courtney/Desktop/c2s2-tape-out-23/openlane/tape_in_mar/runs/23_06_05_15_07/results/signoff/FFTSPIInterconnectRTL.magic.gds
string GDS_START 1901164
<< end >>

