VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO FFTSPIInterconnectRTL
  CLASS BLOCK ;
  FOREIGN FFTSPIInterconnectRTL ;
  ORIGIN 0.000 0.000 ;
  SIZE 1500.000 BY 1500.000 ;
  PIN adapter_parity
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1046.590 0.000 1046.870 4.000 ;
    END
  END adapter_parity
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.130 0.000 747.410 4.000 ;
    END
  END clk
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 975.750 1496.000 976.030 1500.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 785.440 1500.000 786.040 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 472.640 4.000 473.240 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.410 1496.000 824.690 1500.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1497.390 0.000 1497.670 4.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 1496.000 225.770 1500.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1101.640 1500.000 1102.240 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1346.050 0.000 1346.330 4.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1423.330 1496.000 1423.610 1500.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1261.440 1500.000 1262.040 ;
    END
  END io_oeb[18]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.830 1496.000 377.110 1500.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1264.840 4.000 1265.440 ;
    END
  END io_oeb[2]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 312.840 1500.000 313.440 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 788.840 4.000 789.440 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 945.240 1500.000 945.840 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 948.640 4.000 949.240 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1123.870 1496.000 1124.150 1500.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END io_oeb[9]
  PIN master_cs
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.670 0.000 447.950 4.000 ;
    END
  END master_cs
  PIN master_miso
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 1496.000 77.650 1500.000 ;
    END
  END master_miso
  PIN master_mosi
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1197.930 0.000 1198.210 4.000 ;
    END
  END master_mosi
  PIN master_sclk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1275.210 1496.000 1275.490 1500.000 ;
    END
  END master_sclk
  PIN minion_cs
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 153.040 1500.000 153.640 ;
    END
  END minion_cs
  PIN minion_cs_2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END minion_cs_2
  PIN minion_cs_3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 0.000 299.830 4.000 ;
    END
  END minion_cs_3
  PIN minion_miso
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.240 4.000 316.840 ;
    END
  END minion_miso
  PIN minion_miso_2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 469.240 1500.000 469.840 ;
    END
  END minion_miso_2
  PIN minion_miso_3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.010 0.000 599.290 4.000 ;
    END
  END minion_miso_3
  PIN minion_mosi
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1105.040 4.000 1105.640 ;
    END
  END minion_mosi
  PIN minion_mosi_2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1417.840 1500.000 1418.440 ;
    END
  END minion_mosi_2
  PIN minion_mosi_3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.950 1496.000 525.230 1500.000 ;
    END
  END minion_mosi_3
  PIN minion_parity
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.290 1496.000 676.570 1500.000 ;
    END
  END minion_parity
  PIN minion_sclk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 898.470 0.000 898.750 4.000 ;
    END
  END minion_sclk
  PIN minion_sclk_2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 632.440 4.000 633.040 ;
    END
  END minion_sclk_2
  PIN minion_sclk_3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1421.240 4.000 1421.840 ;
    END
  END minion_sclk_3
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 629.040 1500.000 629.640 ;
    END
  END reset
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 1488.080 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 1488.080 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1494.080 1487.925 ;
      LAYER met1 ;
        RECT 0.070 4.460 1497.690 1495.620 ;
      LAYER met2 ;
        RECT 0.100 1495.720 77.090 1496.000 ;
        RECT 77.930 1495.720 225.210 1496.000 ;
        RECT 226.050 1495.720 376.550 1496.000 ;
        RECT 377.390 1495.720 524.670 1496.000 ;
        RECT 525.510 1495.720 676.010 1496.000 ;
        RECT 676.850 1495.720 824.130 1496.000 ;
        RECT 824.970 1495.720 975.470 1496.000 ;
        RECT 976.310 1495.720 1123.590 1496.000 ;
        RECT 1124.430 1495.720 1274.930 1496.000 ;
        RECT 1275.770 1495.720 1423.050 1496.000 ;
        RECT 1423.890 1495.720 1497.660 1496.000 ;
        RECT 0.100 4.280 1497.660 1495.720 ;
        RECT 0.650 3.670 147.930 4.280 ;
        RECT 148.770 3.670 299.270 4.280 ;
        RECT 300.110 3.670 447.390 4.280 ;
        RECT 448.230 3.670 598.730 4.280 ;
        RECT 599.570 3.670 746.850 4.280 ;
        RECT 747.690 3.670 898.190 4.280 ;
        RECT 899.030 3.670 1046.310 4.280 ;
        RECT 1047.150 3.670 1197.650 4.280 ;
        RECT 1198.490 3.670 1345.770 4.280 ;
        RECT 1346.610 3.670 1497.110 4.280 ;
      LAYER met3 ;
        RECT 4.000 1422.240 1496.000 1488.005 ;
        RECT 4.400 1420.840 1496.000 1422.240 ;
        RECT 4.000 1418.840 1496.000 1420.840 ;
        RECT 4.000 1417.440 1495.600 1418.840 ;
        RECT 4.000 1265.840 1496.000 1417.440 ;
        RECT 4.400 1264.440 1496.000 1265.840 ;
        RECT 4.000 1262.440 1496.000 1264.440 ;
        RECT 4.000 1261.040 1495.600 1262.440 ;
        RECT 4.000 1106.040 1496.000 1261.040 ;
        RECT 4.400 1104.640 1496.000 1106.040 ;
        RECT 4.000 1102.640 1496.000 1104.640 ;
        RECT 4.000 1101.240 1495.600 1102.640 ;
        RECT 4.000 949.640 1496.000 1101.240 ;
        RECT 4.400 948.240 1496.000 949.640 ;
        RECT 4.000 946.240 1496.000 948.240 ;
        RECT 4.000 944.840 1495.600 946.240 ;
        RECT 4.000 789.840 1496.000 944.840 ;
        RECT 4.400 788.440 1496.000 789.840 ;
        RECT 4.000 786.440 1496.000 788.440 ;
        RECT 4.000 785.040 1495.600 786.440 ;
        RECT 4.000 633.440 1496.000 785.040 ;
        RECT 4.400 632.040 1496.000 633.440 ;
        RECT 4.000 630.040 1496.000 632.040 ;
        RECT 4.000 628.640 1495.600 630.040 ;
        RECT 4.000 473.640 1496.000 628.640 ;
        RECT 4.400 472.240 1496.000 473.640 ;
        RECT 4.000 470.240 1496.000 472.240 ;
        RECT 4.000 468.840 1495.600 470.240 ;
        RECT 4.000 317.240 1496.000 468.840 ;
        RECT 4.400 315.840 1496.000 317.240 ;
        RECT 4.000 313.840 1496.000 315.840 ;
        RECT 4.000 312.440 1495.600 313.840 ;
        RECT 4.000 157.440 1496.000 312.440 ;
        RECT 4.400 156.040 1496.000 157.440 ;
        RECT 4.000 154.040 1496.000 156.040 ;
        RECT 4.000 152.640 1495.600 154.040 ;
        RECT 4.000 10.715 1496.000 152.640 ;
      LAYER met4 ;
        RECT 498.015 11.735 558.240 1485.625 ;
        RECT 560.640 11.735 635.040 1485.625 ;
        RECT 637.440 11.735 711.840 1485.625 ;
        RECT 714.240 11.735 788.640 1485.625 ;
        RECT 791.040 11.735 865.440 1485.625 ;
        RECT 867.840 11.735 942.240 1485.625 ;
        RECT 944.640 11.735 988.705 1485.625 ;
  END
END FFTSPIInterconnectRTL
END LIBRARY

