VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO FFTSPIInterconnectRTL
  CLASS BLOCK ;
  FOREIGN FFTSPIInterconnectRTL ;
  ORIGIN 0.000 0.000 ;
  SIZE 2320.000 BY 2920.000 ;
  PIN adapter_parity
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2316.000 92.520 2320.000 93.120 ;
    END
  END adapter_parity
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.690 0.000 579.970 4.000 ;
    END
  END clk
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2316.000 274.760 2320.000 275.360 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1610.550 2916.000 1610.830 2920.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1352.950 2916.000 1353.230 2920.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1095.350 2916.000 1095.630 2920.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 837.750 2916.000 838.030 2920.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 580.150 2916.000 580.430 2920.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.550 2916.000 322.830 2920.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.950 2916.000 65.230 2920.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 729.680 4.000 730.280 ;
    END
  END io_oeb[17]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2316.000 639.240 2320.000 639.840 ;
    END
  END io_oeb[1]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2316.000 1003.720 2320.000 1004.320 ;
    END
  END io_oeb[2]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2316.000 1368.200 2320.000 1368.800 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2316.000 1732.680 2320.000 1733.280 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2316.000 2097.160 2320.000 2097.760 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2316.000 2461.640 2320.000 2462.240 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2316.000 2826.120 2320.000 2826.720 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2125.750 2916.000 2126.030 2920.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1868.150 2916.000 1868.430 2920.000 ;
    END
  END io_oeb[9]
  PIN master_cs
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.950 2916.000 709.230 2920.000 ;
    END
  END master_cs
  PIN master_miso
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.350 2916.000 451.630 2920.000 ;
    END
  END master_miso
  PIN master_mosi
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.750 2916.000 194.030 2920.000 ;
    END
  END master_mosi
  PIN master_sclk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2189.640 4.000 2190.240 ;
    END
  END master_sclk
  PIN minion_cs
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2316.000 821.480 2320.000 822.080 ;
    END
  END minion_cs
  PIN minion_cs_2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2316.000 2279.400 2320.000 2280.000 ;
    END
  END minion_cs_2
  PIN minion_cs_3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1739.350 2916.000 1739.630 2920.000 ;
    END
  END minion_cs_3
  PIN minion_miso
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2316.000 1914.920 2320.000 1915.520 ;
    END
  END minion_miso
  PIN minion_miso_2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1996.950 2916.000 1997.230 2920.000 ;
    END
  END minion_miso_2
  PIN minion_miso_3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 966.550 2916.000 966.830 2920.000 ;
    END
  END minion_miso_3
  PIN minion_mosi
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2316.000 1185.960 2320.000 1186.560 ;
    END
  END minion_mosi
  PIN minion_mosi_2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2316.000 2643.880 2320.000 2644.480 ;
    END
  END minion_mosi_2
  PIN minion_mosi_3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1481.750 2916.000 1482.030 2920.000 ;
    END
  END minion_mosi_3
  PIN minion_parity
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2316.000 457.000 2320.000 457.600 ;
    END
  END minion_parity
  PIN minion_sclk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2316.000 1550.440 2320.000 1551.040 ;
    END
  END minion_sclk
  PIN minion_sclk_2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2254.550 2916.000 2254.830 2920.000 ;
    END
  END minion_sclk_2
  PIN minion_sclk_3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1224.150 2916.000 1224.430 2920.000 ;
    END
  END minion_sclk_3
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1739.350 0.000 1739.630 4.000 ;
    END
  END reset
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 2907.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 2907.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 2907.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 2907.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 2907.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 2907.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 2907.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 2907.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 2907.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 2907.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.040 10.640 1558.640 2907.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1710.640 10.640 1712.240 2907.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1864.240 10.640 1865.840 2907.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 2017.840 10.640 2019.440 2907.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 2171.440 10.640 2173.040 2907.920 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 2907.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 2907.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 2907.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 2907.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 2907.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 2907.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 2907.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 2907.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 2907.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 2907.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1633.840 10.640 1635.440 2907.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1787.440 10.640 1789.040 2907.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1941.040 10.640 1942.640 2907.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 2094.640 10.640 2096.240 2907.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 2248.240 10.640 2249.840 2907.920 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 2314.260 2907.765 ;
      LAYER met1 ;
        RECT 4.670 10.640 2315.570 2915.800 ;
      LAYER met2 ;
        RECT 4.690 2915.720 64.670 2916.000 ;
        RECT 65.510 2915.720 193.470 2916.000 ;
        RECT 194.310 2915.720 322.270 2916.000 ;
        RECT 323.110 2915.720 451.070 2916.000 ;
        RECT 451.910 2915.720 579.870 2916.000 ;
        RECT 580.710 2915.720 708.670 2916.000 ;
        RECT 709.510 2915.720 837.470 2916.000 ;
        RECT 838.310 2915.720 966.270 2916.000 ;
        RECT 967.110 2915.720 1095.070 2916.000 ;
        RECT 1095.910 2915.720 1223.870 2916.000 ;
        RECT 1224.710 2915.720 1352.670 2916.000 ;
        RECT 1353.510 2915.720 1481.470 2916.000 ;
        RECT 1482.310 2915.720 1610.270 2916.000 ;
        RECT 1611.110 2915.720 1739.070 2916.000 ;
        RECT 1739.910 2915.720 1867.870 2916.000 ;
        RECT 1868.710 2915.720 1996.670 2916.000 ;
        RECT 1997.510 2915.720 2125.470 2916.000 ;
        RECT 2126.310 2915.720 2254.270 2916.000 ;
        RECT 2255.110 2915.720 2315.550 2916.000 ;
        RECT 4.690 4.280 2315.550 2915.720 ;
        RECT 4.690 4.000 579.410 4.280 ;
        RECT 580.250 4.000 1739.070 4.280 ;
        RECT 1739.910 4.000 2315.550 4.280 ;
      LAYER met3 ;
        RECT 4.000 2827.120 2316.000 2907.845 ;
        RECT 4.000 2825.720 2315.600 2827.120 ;
        RECT 4.000 2644.880 2316.000 2825.720 ;
        RECT 4.000 2643.480 2315.600 2644.880 ;
        RECT 4.000 2462.640 2316.000 2643.480 ;
        RECT 4.000 2461.240 2315.600 2462.640 ;
        RECT 4.000 2280.400 2316.000 2461.240 ;
        RECT 4.000 2279.000 2315.600 2280.400 ;
        RECT 4.000 2190.640 2316.000 2279.000 ;
        RECT 4.400 2189.240 2316.000 2190.640 ;
        RECT 4.000 2098.160 2316.000 2189.240 ;
        RECT 4.000 2096.760 2315.600 2098.160 ;
        RECT 4.000 1915.920 2316.000 2096.760 ;
        RECT 4.000 1914.520 2315.600 1915.920 ;
        RECT 4.000 1733.680 2316.000 1914.520 ;
        RECT 4.000 1732.280 2315.600 1733.680 ;
        RECT 4.000 1551.440 2316.000 1732.280 ;
        RECT 4.000 1550.040 2315.600 1551.440 ;
        RECT 4.000 1369.200 2316.000 1550.040 ;
        RECT 4.000 1367.800 2315.600 1369.200 ;
        RECT 4.000 1186.960 2316.000 1367.800 ;
        RECT 4.000 1185.560 2315.600 1186.960 ;
        RECT 4.000 1004.720 2316.000 1185.560 ;
        RECT 4.000 1003.320 2315.600 1004.720 ;
        RECT 4.000 822.480 2316.000 1003.320 ;
        RECT 4.000 821.080 2315.600 822.480 ;
        RECT 4.000 730.680 2316.000 821.080 ;
        RECT 4.400 729.280 2316.000 730.680 ;
        RECT 4.000 640.240 2316.000 729.280 ;
        RECT 4.000 638.840 2315.600 640.240 ;
        RECT 4.000 458.000 2316.000 638.840 ;
        RECT 4.000 456.600 2315.600 458.000 ;
        RECT 4.000 275.760 2316.000 456.600 ;
        RECT 4.000 274.360 2315.600 275.760 ;
        RECT 4.000 93.520 2316.000 274.360 ;
        RECT 4.000 92.120 2315.600 93.520 ;
        RECT 4.000 10.715 2316.000 92.120 ;
      LAYER met4 ;
        RECT 350.815 24.655 404.640 2906.145 ;
        RECT 407.040 24.655 481.440 2906.145 ;
        RECT 483.840 24.655 558.240 2906.145 ;
        RECT 560.640 24.655 635.040 2906.145 ;
        RECT 637.440 24.655 711.840 2906.145 ;
        RECT 714.240 24.655 788.640 2906.145 ;
        RECT 791.040 24.655 865.440 2906.145 ;
        RECT 867.840 24.655 942.240 2906.145 ;
        RECT 944.640 24.655 1019.040 2906.145 ;
        RECT 1021.440 24.655 1095.840 2906.145 ;
        RECT 1098.240 24.655 1172.640 2906.145 ;
        RECT 1175.040 24.655 1249.440 2906.145 ;
        RECT 1251.840 24.655 1326.240 2906.145 ;
        RECT 1328.640 24.655 1403.040 2906.145 ;
        RECT 1405.440 24.655 1479.840 2906.145 ;
        RECT 1482.240 24.655 1556.640 2906.145 ;
        RECT 1559.040 24.655 1633.440 2906.145 ;
        RECT 1635.840 24.655 1710.240 2906.145 ;
        RECT 1712.640 24.655 1787.040 2906.145 ;
        RECT 1789.440 24.655 1863.840 2906.145 ;
        RECT 1866.240 24.655 1940.640 2906.145 ;
        RECT 1943.040 24.655 2017.440 2906.145 ;
        RECT 2019.840 24.655 2030.145 2906.145 ;
  END
END FFTSPIInterconnectRTL
END LIBRARY

